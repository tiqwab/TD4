module IC74HC32(
    input A,
    input B,
    output wire Y
);

assign Y = A | B;

endmodule
